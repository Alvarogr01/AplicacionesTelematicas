<!DOCTYPE html>
<html lang="es">
    <head>
        <div class="Cursos indra"
            <title>Cursos formativos de Indra </title>
            <link rel="stylesheet" type="text/css" href="Hoja de estilos.css" />
            <meta charset="UTF-8">
        </div>
    </head>
    <body>
        
    
    </body>
</html>
